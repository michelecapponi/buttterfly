LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SWAP IS
	GENERIC( N   : INTEGER:=40);
	PORT (IN_1   : IN SIGNED(N-1 DOWNTO 0);
			IN_2   : IN SIGNED(N-1 DOWNTO 0);
			SW     : IN STD_LOGIC;
			OUT_1  : OUT SIGNED(N-1 DOWNTO 0);
			OUT_2  : OUT SIGNED(N-1 DOWNTO 0));
END SWAP;

ARCHITECTURE BEHAVIOR OF SWAP  IS

BEGIN

PROCESS (IN_1,IN_2,SW)
	BEGIN
		 IF SW = '0' THEN
			 OUT_1<=IN_1;
			 OUT_2<=IN_2;
		ELSE 
			 OUT_1<=IN_2;
			 OUT_2<=IN_1;	
		END IF;
END PROCESS;

END BEHAVIOR;