LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY uROM IS
	PORT(
			ADD : IN STD_LOGIC_VECTOR(3 downto 0);
			ROW : OUT STD_LOGIC_VECTOR(43 downto 0)
		  );
END uROM;

ARCHITECTURE BEHAVIOUR OF uROM IS

BEGIN

PROCESS_OUT : PROCESS(ADD)

BEGIN

CASE ADD IS
	WHEN "0000" => ROW <= "1010000100000000"&"01110"&"0"   &   "1001100100000000"&"00010"&"0";
	WHEN "0001" => ROW <= "1101101100000000"&"00011"&"0"   &   "1111101010000000"&"00100"&"0";
	WHEN "0010" => ROW <= "0001001000000000"&"00101"&"0"   &   "0101001000000000"&"10000"&"1";
	WHEN "0011" => ROW <= "0101011001011000"&"00111"&"0"   &   "0101011001110100"&"01000"&"0";
	WHEN "0100" => ROW <= "0101011000110010"&"01001"&"0"   &   "0101011000110001"&"01110"&"0";
	WHEN "0101" => ROW <= "1001111001011000"&"01011"&"0"   &   "1101101101110100"&"01100"&"0";
	WHEN "0110" => ROW <= "1111101010110010"&"01101"&"0"   &   "0001001000000001"&"00101"&"0";
	WHEN "0111" => ROW <= "1010000100000000"&"01110"&"1"   &   "1011100100000000"&"00001"&"0";
	WHEN "1000" => ROW <= "0101011000110000"&"00110"&"0"   &   "1011111000110000"&"01010"&"0";
	WHEN OTHERS => ROW <= "1010000100000000"&"01110"&"0"   &   "1011100100000000"&"00010"&"0";
END CASE;

END PROCESS;

END BEHAVIOUR;