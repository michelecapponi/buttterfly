LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REG_uAR IS
	PORT (D      : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			CLOCK  : IN STD_LOGIC;
			ENABLE : IN STD_LOGIC;
			RESETN : IN STD_LOGIC;
			Q      : OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END REG_uAR;

ARCHITECTURE BEHAVIOR OF REG_uAR IS

BEGIN
	
	PROCESS (RESETN,CLOCK)
	BEGIN
		 IF RESETN = '0' THEN
			 Q<=(OTHERS=>'0');
		 ELSIF FALLING_EDGE(CLOCK) THEN
			IF (ENABLE = '1') THEN
				Q<=D;
			END IF;
		 END IF;
	END PROCESS;
	
END BEHAVIOR;