LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY LATE_STATUS IS
	PORT(
			CLOCK, RESET_N, START : IN STD_LOGIC;
			SEL_0, SEL_2 : OUT STD_LOGIC_VECTOR(1 downto 0);
			SEL_1, EN_0, EN_7, SHIFT_MULT_N, EN_1, EN_2, SW, SUB_ADD_N, ROUND, EN_3, EN_4, EN_5, EN_6: OUT STD_LOGIC;
			DONE : OUT STD_LOGIC
	);
END LATE_STATUS;

ARCHITECTURE BEHAVIOUR OF LATE_STATUS IS

COMPONENT uROM IS
	PORT(
			ADD : IN STD_LOGIC_VECTOR(3 downto 0);
			ROW : OUT STD_LOGIC_VECTOR(43 downto 0)
		  );
END COMPONENT;

COMPONENT REG_uAR IS
	PORT (D      : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			CLOCK  : IN STD_LOGIC;
			ENABLE : IN STD_LOGIC;
			RESETN : IN STD_LOGIC;
			Q      : OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END COMPONENT;

COMPONENT REG_uIR IS
	PORT (D      : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
			CLOCK  : IN STD_LOGIC;
			ENABLE : IN STD_LOGIC;
			RESETN : IN STD_LOGIC;
			Q      : OUT STD_LOGIC_VECTOR(21 DOWNTO 0));
END COMPONENT;

COMPONENT MUX_2_TO_1_IR is
	GENERIC( N   : INTEGER:=22);
	port(
		  IN_1     : in std_logic_vector(N-1 downto 0);
        IN_2     : in std_logic_vector(N-1 downto 0);
        SEL      : in std_logic;
		  MUX_OUT  : out std_logic_vector(N-1 downto 0));
END COMPONENT;

COMPONENT MUX_2_TO_1_1_BIT is
	port(
		  IN_1     : in std_logic;
        IN_2     : in std_logic;
        SEL      : in std_logic;
		  MUX_OUT  : out std_logic);
end COMPONENT;

SIGNAL MSB_NEXT_ADDRESS, MSB_PRESENT_ADDRESS : STD_LOGIC_VECTOR(3 downto 0);
SIGNAL LSB_NEXT_ADDRESS, LSB_PRESENT_ADDRESS : STD_LOGIC;
SIGNAL uROM_OUT : STD_LOGIC_VECTOR(43 downto 0);
SIGNAL MUX_OUT, uINSTRUCTION, EVEN, ODD : STD_LOGIC_VECTOR(21 downto 0);
SIGNAL CC, LSB_INST_REG : STD_LOGIC;

BEGIN

uAR : REG_uAR PORT MAP(CLOCK=>CLOCK, RESETN=>RESET_N, D(4 downto 1)=>MSB_NEXT_ADDRESS, D(0)=>LSB_NEXT_ADDRESS, ENABLE=>'1', Q(4 downto 1)=>MSB_PRESENT_ADDRESS, Q(0)=>LSB_PRESENT_ADDRESS);

TABLE : uROM PORT MAP (ADD=>MSB_PRESENT_ADDRESS, ROW=>uROM_OUT);

EVEN<=uROM_OUT(43 downto 22);
ODD<=uROM_OUT(21 downto 0);

MUX : MUX_2_TO_1_IR GENERIC MAP (N=>22) PORT MAP(IN_1=>EVEN, IN_2=>ODD, SEL=>LSB_PRESENT_ADDRESS, MUX_OUT=>MUX_OUT);

uIR : REG_uIR PORT MAP(CLOCK=>CLOCK, RESETN=>RESET_N, D=>MUX_OUT, ENABLE=>'1', Q=>uINSTRUCTION);

CC<=uINSTRUCTION(0);
LSB_INST_REG<=uINSTRUCTION(1);
MSB_NEXT_ADDRESS<=uINSTRUCTION(5 downto 2); --dubbio su come vengono messi nella variabile
SEL_0<=uINSTRUCTION(21 downto 20);
SEL_2<=uINSTRUCTION(14 downto 13);
SEL_1<=uINSTRUCTION(19);
EN_0<=uINSTRUCTION(18);
EN_7<=uINSTRUCTION(17);
SHIFT_MULT_N<=uINSTRUCTION(16);
EN_1<=uINSTRUCTION(15);
EN_2<=uINSTRUCTION(15);
SW<=uINSTRUCTION(12);
SUB_ADD_N<=uINSTRUCTION(11);
ROUND<=uINSTRUCTION(10);
EN_3<=uINSTRUCTION(9);
EN_4<=uINSTRUCTION(8);
EN_5<=uINSTRUCTION(7);
EN_6<=uINSTRUCTION(6);
DONE<=uINSTRUCTION(6);

STATUS_PLA : MUX_2_TO_1_1_BIT PORT MAP(IN_2=>START, IN_1=>LSB_INST_REG, SEL=>CC, MUX_OUT=>LSB_NEXT_ADDRESS);

END BEHAVIOUR;